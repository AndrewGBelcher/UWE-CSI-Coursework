module Rom(
	input [3:0]address,
	output logic [23:0]q
);

reg [23:0][7:0]ROM;

always@(address)
begin
	case(address)

		// ones counter
						//bi__ba__ie_we_wa_rae_raa_rbe_rba_alusel_sh_oe__done
		/*4'b0000: q = 25'b001__0001__0_0_00_0_00_0_00_000_00_0__0;
		4'b0001: q = 25'b000__0010__1_1_00_0_00_0_00_000_00_0__0;
		4'b0010: q = 25'b000__0011__0_1_01_1_00_1_00_101_00_0__0;
		4'b0011: q = 25'b000__0100__0_1_10_1_01_0_00_110_00_0__0;
		4'b0100: q = 25'b000__0101__0_1_11_1_00_1_10_001_00_0__0;
		4'b0101: q = 25'b000__0110__0_1_01_1_01_1_11_100_00_0__0;
		4'b0110: q = 25'b010__0100__0_1_00_1_00_0_00_000_10_0__0;
		4'b0111: q = 25'b011__0000__0_0_00_1_01_0_00_000_00_1__1;

		default: q = 25'b001__0001__0_0_00_000_000_000_00_0__0;*/


			//bi__ba__ie_we_wa_rae_raa_rbe_rba_alusel_sh_oe__done
			// 0 pc++ / 1 wait / 2 bnz / 3 reset / 4 b / 5 bn
		4'b0000: q = 24'b001__0001__0_0_00_0_00_0_00_000_00_0__0; // start  		0
		4'b0001: q = 24'b000__0010__1_1_00_0_00_0_00_000_00_0__0; // load a		1
		4'b0010: q = 24'b000__0011__1_1_01_0_00_0_00_000_00_0__0; // load b		2
			
		4'b0011: q = 24'b010__0101__0_1_10_1_00_1_01_101_00_0__0; // a - b = c		3
		4'b0100: q = 24'b001__0000__0_0_00_1_00_0_00_000_00_1__1; // done s4		4
		4'b0101: q = 24'b101__0111__0_0_00_1_10_0_00_000_00_0__0; // is neg? aka a < b	5

		4'b0110: q = 24'b100__0011__0_1_00_1_10_0_00_000_00_0__0; // a > b a = c	6

		4'b0111: q = 24'b000__1000__0_1_11_1_00_0_00_000_00_0__0; // d = a		7
		4'b1000: q = 24'b000__1001__0_1_00_1_01_0_00_000_00_0__0; // a = b		8
		4'b1001: q = 24'b100__0011__0_1_01_1_11_0_00_000_00_0__0; // b = d goto s3	9

	endcase
end
endmodule