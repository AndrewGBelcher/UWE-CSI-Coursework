//module alu (input alu_1,
//				input alu_2,
//				input alu_3