//module gcd_controller(input clk,
//							 input reset,
//							 input start,
//							 input done
//							 );
//				
//
//				
//endmodule;